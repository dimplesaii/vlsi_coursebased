module dadda_16(output [31:0]y, input [15:0]a,b);
wire [14:0] hs,hc;
wire [194:0] fs,fc;
wire [255:0]p;
wire [30:1]c;
genvar i,j;
generate
for(i=0; i<16; i=i+1) begin: pr
	for(j=0; j<16; j=j+1)begin:pc
		assign p[i+(j*16)] = a[i] & b[j]; 		//Partial Product Generation
	end
end
endgenerate
	
//Reduction Stage 1: Dj = 13
HA h0 (hs[0], hc[0], p[13], p[28]);	
FA f0 (fs[0], fc[0], hc[0], p[14], p[29]);
HA h1 (hs[1], hc[1], p[44], p[59]);
FA f1 (fs[1], fc[1], hc[1], fc[0], p[15]);
FA f2 (fs[2], fc[2], p[30], p[45], p[60]);
HA h2 (hs[2], hc[2], p[75], p[90]);
FA f3 (fs[3], fc[3], hc[2], fc[2], fc[1]);
FA f4 (fs[4], fc[4], p[31], p[46], p[61]);
HA h3 (hs[3], hc[3], p[76], p[91]);
FA f5 (fs[5], fc[5], hc[3], fc[4], fc[3]);
FA f6 (fs[6], fc[6], p[47], p[62], p[77]);
FA f7 (fs[7], fc[7], fc[6], fc[5], p[63]);
	
//Reduction Stage 2: Dj = 9
HA h4 (hs[4], hc[4], p[9], p[24]);
FA f8 (fs[8], fc[8], hc[4], p[10], p[25]);
HA h5 (hs[5], hc[5], p[40], p[55]);
FA f9 (fs[9], fc[9], hc[5], fc[8], p[11]);
FA f10 (fs[10], fc[10], p[26], p[41], p[56]);
HA h6 (hs[6], hc[6], p[71], p[86]);
FA f11 (fs[11], fc[11], hc[6], fc[10], fc[9]);
FA f12 (fs[12], fc[12], p[12], p[27], p[42]);
FA f13 (fs[13], fc[13], p[57], p[72], p[87]);
HA h7 (hs[7], hc[7], p[102], p[117]);
FA f14 (fs[14], fc[14], hc[7], fc[13], fc[12]);
FA f15 (fs[15], fc[15], fc[11], hs[0], p[43]);
FA f16 (fs[16], fc[16], p[58], p[73], p[88]);
FA f17 (fs[17], fc[17], p[103], p[118], p[133]);
FA f18 (fs[18], fc[18], fc[17], fc[16], fc[15]);
FA f19 (fs[19], fc[19], fc[14], fs[0], hs[1]);
FA f20 (fs[20], fc[20], p[74], p[89], p[104]);
FA f21 (fs[21], fc[21], p[119], p[134], p[149]);
FA f22 (fs[22], fc[22], fc[21], fc[20], fc[19]);
FA f23 (fs[23], fc[23], fc[18], fs[2], fs[1]);
FA f24 (fs[24], fc[24], hs[2], p[105], p[120]);
FA f25 (fs[25], fc[25], p[135], p[150], p[165]);
FA f26 (fs[26], fc[26], fc[25], fc[24], fc[23]);
FA f27 (fs[27], fc[27], fc[22], fs[4], fs[3]);
FA f28 (fs[28], fc[28], hs[3], p[106], p[121]);
FA f29 (fs[29], fc[29], p[136], p[151], p[166]);
FA f30 (fs[30], fc[30], fc[29], fc[28], fc[27]);
FA f31 (fs[31], fc[31], fc[26], fs[6], fs[5]);
FA f32 (fs[32], fc[32], p[92], p[107], p[122]);
FA f33 (fs[33], fc[33], p[137], p[152], p[167]);
FA f34 (fs[34], fc[34], fc[33], fc[32], fc[31]);
FA f35 (fs[35], fc[35], fc[30], fs[7], p[78]);
FA f36 (fs[36], fc[36], p[93], p[108], p[123]);
FA f37 (fs[37], fc[37], p[138], p[153], p[168]);
FA f38 (fs[38], fc[38], fc[37], fc[36], fc[35]);
FA f39 (fs[39], fc[39], fc[34], fc[7], p[79]);
FA f40 (fs[40], fc[40], p[94], p[109], p[124]);
FA f41 (fs[41], fc[41], p[139], p[154], p[169]);
FA f42 (fs[42], fc[42], fc[41], fc[40], fc[39]);
FA f43 (fs[43], fc[43], fc[38], p[95], p[110]);
FA f44 (fs[44], fc[44], p[125], p[140], p[155]);
FA f45 (fs[45], fc[45], fc[44], fc[43], fc[42]);
FA f46 (fs[46], fc[46], p[111], p[126], p[141]);
FA f47 (fs[47], fc[47], fc[46], fc[45], p[127]);
	
//Reduction Stage 3: Dj = 6
HA h8 (hs[8], hc[8], p[6], p[21]);
FA f48 (fs[48], fc[48], hc[8], p[7], p[22]);
HA h9 (hs[9], hc[9], p[37], p[52]);
FA f49 (fs[49], fc[49], hc[9], fc[48], p[8]);
FA f50 (fs[50], fc[50], p[23], p[38], p[53]);
HA h10 (hs[10], hc[10], p[68], p[83]);
FA f51 (fs[51], fc[51], hc[10], fc[50], fc[49]);
FA f52 (fs[52], fc[52], hs[4], p[39], p[54]);
FA f53 (fs[53], fc[53], p[69], p[84], p[99]);
FA f54 (fs[54], fc[54], fc[53], fc[52], fc[51]);
FA f55 (fs[55], fc[55], fs[8], hs[5], p[70]);
FA f56 (fs[56], fc[56], p[85], p[100], p[115]);
FA f57 (fs[57], fc[57], fc[56], fc[55], fc[54]);
FA f58 (fs[58], fc[58], fs[9], fs[10], hs[6]);
FA f59 (fs[59], fc[59], p[101], p[116], p[131]);
FA f60 (fs[60], fc[60], fc[59], fc[58], fc[57]);
FA f61 (fs[61], fc[61], fs[11], fs[12], fs[13]);
FA f62 (fs[62], fc[62], hs[7], p[132], p[147]);
FA f63 (fs[63], fc[63], fc[62], fc[61], fc[60]);
FA f64 (fs[64], fc[64], fs[14], fs[15], fs[16]);
FA f65 (fs[65], fc[65], fs[17], p[148], p[163]);
FA f66 (fs[66], fc[66], fc[65], fc[64], fc[63]);
FA f67 (fs[67], fc[67], fs[18], fs[19], fs[20]);
FA f68 (fs[68], fc[68], fs[21], p[164], p[179]);
FA f69 (fs[69], fc[69], fc[68], fc[67], fc[66]);
FA f70 (fs[70], fc[70], fs[22], fs[23], fs[24]);
FA f71 (fs[71], fc[71], fs[25], p[180], p[195]);
FA f72 (fs[72], fc[72], fc[71], fc[70], fc[69]);
FA f73 (fs[73], fc[73], fs[26], fs[27], fs[28]);
FA f74 (fs[74], fc[74], fs[29], p[181], p[196]);
FA f75 (fs[75], fc[75], fc[74], fc[73], fc[72]);
FA f76 (fs[76], fc[76], fs[30], fs[31], fs[32]);
FA f77 (fs[77], fc[77], fs[33], p[182], p[197]);
FA f78 (fs[78], fc[78], fc[77], fc[76], fc[75]);
FA f79 (fs[79], fc[79], fs[34], fs[35], fs[36]);
FA f80 (fs[80], fc[80], fs[37], p[183], p[198]);
FA f81 (fs[81], fc[81], fc[80], fc[79], fc[78]);
FA f82 (fs[82], fc[82], fs[38], fs[39], fs[40]);
FA f83 (fs[83], fc[83], fs[41], p[184], p[199]);
FA f84 (fs[84], fc[84], fc[83], fc[82], fc[81]);
FA f85 (fs[85], fc[85], fs[42], fs[43], fs[44]);
FA f86 (fs[86], fc[86], p[170], p[185], p[200]);
FA f87 (fs[87], fc[87], fc[86], fc[85], fc[84]);
FA f88 (fs[88], fc[88], fs[45], fs[46], p[156]);
FA f89 (fs[89], fc[89], p[171], p[186], p[201]);
FA f90 (fs[90], fc[90], fc[89], fc[88], fc[87]);
FA f91 (fs[91], fc[91], fs[47], p[142], p[157]);
FA f92 (fs[92], fc[92], p[172], p[187], p[202]);
FA f93 (fs[93], fc[93], fc[92], fc[91], fc[90]);
FA f94 (fs[94], fc[94], fc[47], p[143], p[158]);
FA f95 (fs[95], fc[95], p[173], p[188], p[203]);
FA f96 (fs[96], fc[96], fc[95], fc[94], fc[93]);
FA f97 (fs[97], fc[97], p[159], p[174], p[189]);
FA f98 (fs[98], fc[98], fc[97], fc[96], fc[175]);
	
//Reduction Stage 4: Dj = 4
HA h11 (hs[11], hc[11], p[4], p[19]);
FA f99 (fs[99], fc[99], hc[11], p[5], p[20]);
HA h12 (hs[12], hc[12], p[35], p[50]);
FA f100 (fs[100], fc[100], hc[12], fc[99], hs[8]);
FA f101 (fs[101], fc[101], p[36], p[51], p[66]);
FA f102 (fs[102], fc[102], fc[101], fc[100], fs[48]);
FA f103 (fs[103], fc[103], hs[9], p[67], p[82]);
FA f104 (fs[104], fc[104], fc[103], fc[102], fs[49]);
FA f105 (fs[105], fc[105], fs[50], hs[10], p[98]);
FA f106 (fs[106], fc[106], fc[105], fc[104], fs[51]);
FA f107 (fs[107], fc[107], fs[52], fs[53], p[114]);
FA f108 (fs[108], fc[108], fc[107], fc[106], fs[54]);
FA f109 (fs[109], fc[109], fs[55], fs[56], p[130]);
FA f110 (fs[110], fc[110], fc[109], fc[108], fs[57]);
FA f111 (fs[111], fc[111], fs[58], fs[59], p[146]);
FA f112 (fs[112], fc[112], fc[111], fc[110], fs[60]);
FA f113 (fs[113], fc[113], fs[61], fs[62], p[162]);
FA f114 (fs[114], fc[114], fc[113], fc[112], fs[63]);
FA f115 (fs[115], fc[115], fs[64], fs[65], p[178]);
FA f116 (fs[116], fc[116], fc[115], fc[114], fs[66]);
FA f117 (fs[117], fc[117], fs[67], fs[68], p[194]);
FA f118 (fs[118], fc[118], fc[117], fc[116], fs[69]);
FA f119 (fs[119], fc[119], fs[70], fs[71], p[210]);
FA f120 (fs[120], fc[120], fc[119], fc[118], fs[72]);
FA f121 (fs[121], fc[121], fs[73], fs[74], p[211]);
FA f122 (fs[122], fc[122], fc[121], fc[120], fs[75]);
FA f123 (fs[123], fc[123], fs[76], fs[77], p[212]);
FA f124 (fs[124], fc[124], fc[123], fc[122], fs[78]);
FA f125 (fs[125], fc[125], fs[79], fs[80], p[213]);
FA f126 (fs[126], fc[126], fc[125], fc[124], fs[81]);
FA f127 (fs[127], fc[127], fs[82], fs[83], p[214]);
FA f128 (fs[128], fc[128], fc[127], fc[126], fs[84]);
FA f129 (fs[129], fc[129], fs[85], fs[86], p[215]);
FA f130 (fs[130], fc[130], fc[129], fc[128], fs[87]);
FA f131 (fs[131], fc[131], fs[88], fs[89], p[216]);
FA f132 (fs[132], fc[132], fc[131], fc[130], fs[90]);
FA f133 (fs[133], fc[133], fs[91], fs[92], p[217]);
FA f134 (fs[134], fc[134], fc[133], fc[132], fs[93]);
FA f135 (fs[135], fc[135], fs[94], fs[95], p[218]);
FA f136 (fs[136], fc[136], fc[135], fc[134], fs[96]);
FA f137 (fs[137], fc[137], fs[97], p[204], p[219]);
FA f138 (fs[138], fc[138], fc[137], fc[136], fs[98]);
FA f139 (fs[139], fc[139], p[190], p[205], p[220]);
FA f140 (fs[140], fc[140], fc[139], fc[138], fc[98]);
FA f141 (fs[141], fc[141], p[191], p[206], p[221]);
FA f142 (fs[142], fc[142], fc[141], fc[140], p[207]);
	
//Reduction Stage 5: Dj = 3
HA h13 (hs[13], hc[13], p[3], p[18]);
FA f143 (fs[143], fc[143], hc[13], hs[11], p[34]);
FA f144 (fs[144], fc[144], fc[143], fs[99], hs[12]);
FA f145 (fs[145], fc[145], fc[144], fs[101], fs[100]);
FA f146 (fs[146], fc[146], fc[145], fs[103], fs[102]);
FA f147 (fs[147], fc[147], fc[146], fs[105], fs[104]);
FA f148 (fs[148], fc[148], fc[147], fs[107], fs[106]);
FA f149 (fs[149], fc[149], fc[148], fs[109], fs[108]);
FA f150 (fs[150], fc[150], fc[149], fs[111], fs[110]);
FA f151 (fs[151], fc[151], fc[150], fs[113], fs[112]);
FA f152 (fs[152], fc[152], fc[151], fs[115], fs[114]);
FA f153 (fs[153], fc[153], fc[152], fs[117], fs[116]);
FA f154 (fs[154], fc[154], fc[153], fs[119], fs[118]);
FA f155 (fs[155], fc[155], fc[154], fs[121], fs[120]);
FA f156 (fs[156], fc[156], fc[155], fs[123], fs[122]);
FA f157 (fs[157], fc[157], fc[156], fs[125], fs[124]);
FA f158 (fs[158], fc[158], fc[157], fs[127], fs[126]);
FA f159 (fs[159], fc[159], fc[158], fs[129], fs[128]);
FA f160 (fs[160], fc[160], fc[159], fs[131], fs[130]);
FA f161 (fs[161], fc[161], fc[160], fs[133], fs[132]);
FA f162 (fs[162], fc[162], fc[161], fs[135], fs[134]);
FA f163 (fs[163], fc[163], fc[162], fs[137], fs[136]);
FA f164 (fs[164], fc[164], fc[163], fs[139], fs[138]);
FA f165 (fs[165], fc[165], fc[164], fs[141], fs[140]);
FA f166 (fs[166], fc[166], fc[165], fs[142], p[222]);
FA f167 (fs[167], fc[167], fc[166], fc[142], p[223]);
	
//Reduction Stage 6: Dj = 2
HA h14 (hs[14], hc[14], p[2], p[17]);
FA f168 (fs[168], fc[168], hc[14], hs[13], p[33]);
FA f169 (fs[169], fc[169], fc[168], fs[143], p[49]);
FA f170 (fs[170], fc[170], fc[169], fs[144], p[65]);
FA f171 (fs[171], fc[171], fc[170], fs[145], p[81]);
FA f172 (fs[172], fc[172], fc[171], fs[146], p[97]);
FA f173 (fs[173], fc[173], fc[172], fs[147], p[113]);
FA f174 (fs[174], fc[174], fc[173], fs[148], p[129]);
FA f175 (fs[175], fc[175], fc[174], fs[149], p[145]);
FA f176 (fs[176], fc[176], fc[175], fs[150], p[161]);
FA f177 (fs[177], fc[177], fc[176], fs[151], p[177]);
FA f178 (fs[178], fc[178], fc[177], fs[152], p[193]);
FA f179 (fs[179], fc[179], fc[178], fs[153], p[209]);
FA f180 (fs[180], fc[180], fc[179], fs[154], p[225]);
FA f181 (fs[181], fc[181], fc[180], fs[155], p[226]);
FA f182 (fs[182], fc[182], fc[181], fs[156], p[227]);
FA f183 (fs[183], fc[183], fc[182], fs[157], p[228]);
FA f184 (fs[184], fc[184], fc[183], fs[158], p[229]);
FA f185 (fs[185], fc[185], fc[184], fs[159], p[230]);
FA f186 (fs[186], fc[186], fc[185], fs[160], p[231]);
FA f187 (fs[187], fc[187], fc[186], fs[161], p[232]);
FA f188 (fs[188], fc[188], fc[187], fs[162], p[233]);
FA f189 (fs[189], fc[189], fc[188], fs[163], p[234]);
FA f190 (fs[190], fc[190], fc[189], fs[164], p[235]);
FA f191 (fs[191], fc[191], fc[190], fs[165], p[236]);
FA f192 (fs[192], fc[192], fc[191], fs[166], p[237]);
FA f193 (fs[193], fc[193], fc[192], fs[167], p[238]);
FA f194 (fs[194], fc[194], fc[193], fs[167], p[239]);
	
//Output Vector Generation
buf r0  (y[0], p[0]);
FA  r1  (y[1], c[1], p[1], p[16], 1'b0);
FA  r2  (y[2], c[2], hs[14], p[32], c[1]);
FA  r3  (y[3], c[3], fs[168], p[48], c[2]);
FA  r4  (y[4], c[4], fs[169], p[64], c[3]);
FA  r5  (y[5], c[5], fs[170], p[80], c[4]);
FA  r6  (y[6], c[6], fs[171], p[96], c[5]);
FA  r7  (y[7], c[7], fs[172], p[112], c[6]);
FA  r8  (y[8], c[8], fs[173], p[128], c[7]);
FA  r9  (y[9], c[9], fs[174], p[144], c[8]);
FA  r10 (y[10], c[10], fs[175], p[160], c[9]);
FA  r11 (y[11], c[11], fs[176], p[176], c[10]);
FA  r12 (y[12], c[12], fs[177], p[192], c[11]);
FA  r13 (y[13], c[13], fs[178], p[208], c[12]);
FA  r14 (y[14], c[14], fs[179], p[224], c[13]);
FA  r15 (y[15], c[15], fs[180], p[240], c[14]);
FA  r16 (y[16], c[16], fs[181], p[241], c[15]);
FA  r17 (y[17], c[17], fs[182], p[242], c[16]);
FA  r18 (y[18], c[18], fs[183], p[243], c[17]);
FA  r19 (y[19], c[19], fs[184], p[244], c[18]);
FA  r20 (y[20], c[20], fs[185], p[245], c[19]);
FA  r21 (y[21], c[21], fs[186], p[246], c[20]);
FA  r22 (y[22], c[22], fs[187], p[247], c[21]);
FA  r23 (y[23], c[23], fs[188], p[248], c[22]);
FA  r24 (y[24], c[24], fs[189], p[249], c[23]);
FA  r25 (y[25], c[25], fs[190], p[250], c[24]);
FA  r26 (y[26], c[26], fs[191], p[251], c[25]);
FA  r27 (y[27], c[27], fs[192], p[252], c[26]);
FA  r28 (y[28], c[28], fs[193], p[253], c[27]);
FA  r29 (y[29], c[29], fs[194], p[254], c[28]);
FA  r30 (y[30], c[30], fc[194], p[255], c[29]);
buf r31 (y[31], c[30]);
endmodule

//Full Adder Module
module FA (output s, co, input a, b, ci);
assign s=a^b^ci;
assign co=(a&b)|(b&ci)|(ci&a);
endmodule 

//Half Adder Module
module HA (output s, c, input a, b);
assign s=a^b;
assign c=a&b;
endmodule 
